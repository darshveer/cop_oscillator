* Auto-testbench (planar graph mapped to RO grid)

.include "ptm_45nm_lp.l"
.include "inv.subckt"
.include "nand.subckt"
.include "ring_osc.subckt"
.include "coupling.subckt"
.include "myfile.cir"

Xdut EN_RO_0_0 EN_RO_0_1 EN_RO_0_2 EN_RO_0_3 EN_RO_0_4 EN_RO_0_5 EN_RO_0_6 EN_RO_0_7 EN_RO_0_8 EN_RO_0_9 EN_RO_1_0 EN_RO_1_1 EN_RO_1_2 EN_RO_1_3 EN_RO_1_4 EN_RO_1_5 EN_RO_1_6 EN_RO_1_7 EN_RO_1_8 EN_RO_1_9 EN_RO_2_0 EN_RO_2_1 EN_RO_2_2 EN_RO_2_3 EN_RO_2_4 EN_RO_2_5 EN_RO_2_6 EN_RO_2_7 EN_RO_2_8 EN_RO_2_9 EN_RO_3_0 EN_RO_3_1 EN_RO_3_2 EN_RO_3_3 EN_RO_3_4 EN_RO_3_5 EN_RO_3_6 EN_RO_3_7 EN_RO_3_8 EN_RO_3_9 EN_RO_4_0 EN_RO_4_1 EN_RO_4_2 EN_RO_4_3 EN_RO_4_4 EN_RO_4_5 EN_RO_4_6 EN_RO_4_7 EN_RO_4_8 EN_RO_4_9 EN_RO_5_0 EN_RO_5_1 EN_RO_5_2 EN_RO_5_3 EN_RO_5_4 EN_RO_5_5 EN_RO_5_6 EN_RO_5_7 EN_RO_5_8 EN_RO_5_9 EN_RO_6_0 EN_RO_6_1 EN_RO_6_2 EN_RO_6_3 EN_RO_6_4 EN_RO_6_5 EN_RO_6_6 EN_RO_6_7 EN_RO_6_8 EN_RO_6_9 EN_RO_7_0 EN_RO_7_1 EN_RO_7_2 EN_RO_7_3 EN_RO_7_4 EN_RO_7_5 EN_RO_7_6 EN_RO_7_7 EN_RO_7_8 EN_RO_7_9 EN_RO_8_0 EN_RO_8_1 EN_RO_8_2 EN_RO_8_3 EN_RO_8_4 EN_RO_8_5 EN_RO_8_6 EN_RO_8_7 EN_RO_8_8 EN_RO_8_9 EN_RO_9_0 EN_RO_9_1 EN_RO_9_2 EN_RO_9_3 EN_RO_9_4 EN_RO_9_5 EN_RO_9_6 EN_RO_9_7 EN_RO_9_8 EN_RO_9_9 EN_C_0_0__0_1 EN_C_0_0__1_0 EN_C_0_1__0_2 EN_C_0_1__1_0 EN_C_0_1__1_1 EN_C_0_2__0_3 EN_C_0_2__1_1 EN_C_0_2__1_2 EN_C_0_3__0_4 EN_C_0_3__1_2 EN_C_0_3__1_3 EN_C_0_4__0_5 EN_C_0_4__1_3 EN_C_0_4__1_4 EN_C_0_5__0_6 EN_C_0_5__1_4 EN_C_0_5__1_5 EN_C_0_6__0_7 EN_C_0_6__1_5 EN_C_0_6__1_6 EN_C_0_7__0_8 EN_C_0_7__1_6 EN_C_0_7__1_7 EN_C_0_8__0_9 EN_C_0_8__1_7 EN_C_0_8__1_8 EN_C_0_9__1_8 EN_C_0_9__1_9 EN_C_1_0__1_1 EN_C_1_0__2_0 EN_C_1_0__2_1 EN_C_1_1__1_2 EN_C_1_1__2_1 EN_C_1_1__2_2 EN_C_1_2__1_3 EN_C_1_2__2_2 EN_C_1_2__2_3 EN_C_1_3__1_4 EN_C_1_3__2_3 EN_C_1_3__2_4 EN_C_1_4__1_5 EN_C_1_4__2_4 EN_C_1_4__2_5 EN_C_1_5__1_6 EN_C_1_5__2_5 EN_C_1_5__2_6 EN_C_1_6__1_7 EN_C_1_6__2_6 EN_C_1_6__2_7 EN_C_1_7__1_8 EN_C_1_7__2_7 EN_C_1_7__2_8 EN_C_1_8__1_9 EN_C_1_8__2_8 EN_C_1_8__2_9 EN_C_1_9__2_9 EN_C_2_0__2_1 EN_C_2_0__3_0 EN_C_2_1__2_2 EN_C_2_1__3_0 EN_C_2_1__3_1 EN_C_2_2__2_3 EN_C_2_2__3_1 EN_C_2_2__3_2 EN_C_2_3__2_4 EN_C_2_3__3_2 EN_C_2_3__3_3 EN_C_2_4__2_5 EN_C_2_4__3_3 EN_C_2_4__3_4 EN_C_2_5__2_6 EN_C_2_5__3_4 EN_C_2_5__3_5 EN_C_2_6__2_7 EN_C_2_6__3_5 EN_C_2_6__3_6 EN_C_2_7__2_8 EN_C_2_7__3_6 EN_C_2_7__3_7 EN_C_2_8__2_9 EN_C_2_8__3_7 EN_C_2_8__3_8 EN_C_2_9__3_8 EN_C_2_9__3_9 EN_C_3_0__3_1 EN_C_3_0__4_0 EN_C_3_0__4_1 EN_C_3_1__3_2 EN_C_3_1__4_1 EN_C_3_1__4_2 EN_C_3_2__3_3 EN_C_3_2__4_2 EN_C_3_2__4_3 EN_C_3_3__3_4 EN_C_3_3__4_3 EN_C_3_3__4_4 EN_C_3_4__3_5 EN_C_3_4__4_4 EN_C_3_4__4_5 EN_C_3_5__3_6 EN_C_3_5__4_5 EN_C_3_5__4_6 EN_C_3_6__3_7 EN_C_3_6__4_6 EN_C_3_6__4_7 EN_C_3_7__3_8 EN_C_3_7__4_7 EN_C_3_7__4_8 EN_C_3_8__3_9 EN_C_3_8__4_8 EN_C_3_8__4_9 EN_C_3_9__4_9 EN_C_4_0__4_1 EN_C_4_0__5_0 EN_C_4_1__4_2 EN_C_4_1__5_0 EN_C_4_1__5_1 EN_C_4_2__4_3 EN_C_4_2__5_1 EN_C_4_2__5_2 EN_C_4_3__4_4 EN_C_4_3__5_2 EN_C_4_3__5_3 EN_C_4_4__4_5 EN_C_4_4__5_3 EN_C_4_4__5_4 EN_C_4_5__4_6 EN_C_4_5__5_4 EN_C_4_5__5_5 EN_C_4_6__4_7 EN_C_4_6__5_5 EN_C_4_6__5_6 EN_C_4_7__4_8 EN_C_4_7__5_6 EN_C_4_7__5_7 EN_C_4_8__4_9 EN_C_4_8__5_7 EN_C_4_8__5_8 EN_C_4_9__5_8 EN_C_4_9__5_9 EN_C_5_0__5_1 EN_C_5_0__6_0 EN_C_5_0__6_1 EN_C_5_1__5_2 EN_C_5_1__6_1 EN_C_5_1__6_2 EN_C_5_2__5_3 EN_C_5_2__6_2 EN_C_5_2__6_3 EN_C_5_3__5_4 EN_C_5_3__6_3 EN_C_5_3__6_4 EN_C_5_4__5_5 EN_C_5_4__6_4 EN_C_5_4__6_5 EN_C_5_5__5_6 EN_C_5_5__6_5 EN_C_5_5__6_6 EN_C_5_6__5_7 EN_C_5_6__6_6 EN_C_5_6__6_7 EN_C_5_7__5_8 EN_C_5_7__6_7 EN_C_5_7__6_8 EN_C_5_8__5_9 EN_C_5_8__6_8 EN_C_5_8__6_9 EN_C_5_9__6_9 EN_C_6_0__6_1 EN_C_6_0__7_0 EN_C_6_1__6_2 EN_C_6_1__7_0 EN_C_6_1__7_1 EN_C_6_2__6_3 EN_C_6_2__7_1 EN_C_6_2__7_2 EN_C_6_3__6_4 EN_C_6_3__7_2 EN_C_6_3__7_3 EN_C_6_4__6_5 EN_C_6_4__7_3 EN_C_6_4__7_4 EN_C_6_5__6_6 EN_C_6_5__7_4 EN_C_6_5__7_5 EN_C_6_6__6_7 EN_C_6_6__7_5 EN_C_6_6__7_6 EN_C_6_7__6_8 EN_C_6_7__7_6 EN_C_6_7__7_7 EN_C_6_8__6_9 EN_C_6_8__7_7 EN_C_6_8__7_8 EN_C_6_9__7_8 EN_C_6_9__7_9 EN_C_7_0__7_1 EN_C_7_0__8_0 EN_C_7_0__8_1 EN_C_7_1__7_2 EN_C_7_1__8_1 EN_C_7_1__8_2 EN_C_7_2__7_3 EN_C_7_2__8_2 EN_C_7_2__8_3 EN_C_7_3__7_4 EN_C_7_3__8_3 EN_C_7_3__8_4 EN_C_7_4__7_5 EN_C_7_4__8_4 EN_C_7_4__8_5 EN_C_7_5__7_6 EN_C_7_5__8_5 EN_C_7_5__8_6 EN_C_7_6__7_7 EN_C_7_6__8_6 EN_C_7_6__8_7 EN_C_7_7__7_8 EN_C_7_7__8_7 EN_C_7_7__8_8 EN_C_7_8__7_9 EN_C_7_8__8_8 EN_C_7_8__8_9 EN_C_7_9__8_9 EN_C_8_0__8_1 EN_C_8_0__9_0 EN_C_8_1__8_2 EN_C_8_1__9_0 EN_C_8_1__9_1 EN_C_8_2__8_3 EN_C_8_2__9_1 EN_C_8_2__9_2 EN_C_8_3__8_4 EN_C_8_3__9_2 EN_C_8_3__9_3 EN_C_8_4__8_5 EN_C_8_4__9_3 EN_C_8_4__9_4 EN_C_8_5__8_6 EN_C_8_5__9_4 EN_C_8_5__9_5 EN_C_8_6__8_7 EN_C_8_6__9_5 EN_C_8_6__9_6 EN_C_8_7__8_8 EN_C_8_7__9_6 EN_C_8_7__9_7 EN_C_8_8__8_9 EN_C_8_8__9_7 EN_C_8_8__9_8 EN_C_8_9__9_8 EN_C_8_9__9_9 EN_C_9_0__9_1 EN_C_9_1__9_2 EN_C_9_2__9_3 EN_C_9_3__9_4 EN_C_9_4__9_5 EN_C_9_5__9_6 EN_C_9_6__9_7 EN_C_9_7__9_8 EN_C_9_8__9_9 N_0_0_1 N_0_1_1 N_0_2_1 N_0_3_1 N_0_4_1 N_0_5_1 N_0_6_1 N_0_7_1 N_0_8_1 N_0_9_1 N_1_0_1 N_1_1_1 N_1_2_1 N_1_3_1 N_1_4_1 N_1_5_1 N_1_6_1 N_1_7_1 N_1_8_1 N_1_9_1 N_2_0_1 N_2_1_1 N_2_2_1 N_2_3_1 N_2_4_1 N_2_5_1 N_2_6_1 N_2_7_1 N_2_8_1 N_2_9_1 N_3_0_1 N_3_1_1 N_3_2_1 N_3_3_1 N_3_4_1 N_3_5_1 N_3_6_1 N_3_7_1 N_3_8_1 N_3_9_1 N_4_0_1 N_4_1_1 N_4_2_1 N_4_3_1 N_4_4_1 N_4_5_1 N_4_6_1 N_4_7_1 N_4_8_1 N_4_9_1 N_5_0_1 N_5_1_1 N_5_2_1 N_5_3_1 N_5_4_1 N_5_5_1 N_5_6_1 N_5_7_1 N_5_8_1 N_5_9_1 N_6_0_1 N_6_1_1 N_6_2_1 N_6_3_1 N_6_4_1 N_6_5_1 N_6_6_1 N_6_7_1 N_6_8_1 N_6_9_1 N_7_0_1 N_7_1_1 N_7_2_1 N_7_3_1 N_7_4_1 N_7_5_1 N_7_6_1 N_7_7_1 N_7_8_1 N_7_9_1 N_8_0_1 N_8_1_1 N_8_2_1 N_8_3_1 N_8_4_1 N_8_5_1 N_8_6_1 N_8_7_1 N_8_8_1 N_8_9_1 N_9_0_1 N_9_1_1 N_9_2_1 N_9_3_1 N_9_4_1 N_9_5_1 N_9_6_1 N_9_7_1 N_9_8_1 N_9_9_1 vdd gnd RING_OSC_NETWORK

* RO enables
V_EN_RO_0_0 EN_RO_0_0 gnd 1
V_EN_RO_0_1 EN_RO_0_1 gnd 0
V_EN_RO_0_2 EN_RO_0_2 gnd 1
V_EN_RO_0_3 EN_RO_0_3 gnd 0
V_EN_RO_0_4 EN_RO_0_4 gnd 0
V_EN_RO_0_5 EN_RO_0_5 gnd 0
V_EN_RO_0_6 EN_RO_0_6 gnd 0
V_EN_RO_0_7 EN_RO_0_7 gnd 1
V_EN_RO_0_8 EN_RO_0_8 gnd 1
V_EN_RO_0_9 EN_RO_0_9 gnd 0
V_EN_RO_1_0 EN_RO_1_0 gnd 1
V_EN_RO_1_1 EN_RO_1_1 gnd 0
V_EN_RO_1_2 EN_RO_1_2 gnd 0
V_EN_RO_1_3 EN_RO_1_3 gnd 1
V_EN_RO_1_4 EN_RO_1_4 gnd 1
V_EN_RO_1_5 EN_RO_1_5 gnd 1
V_EN_RO_1_6 EN_RO_1_6 gnd 0
V_EN_RO_1_7 EN_RO_1_7 gnd 0
V_EN_RO_1_8 EN_RO_1_8 gnd 0
V_EN_RO_1_9 EN_RO_1_9 gnd 0
V_EN_RO_2_0 EN_RO_2_0 gnd 1
V_EN_RO_2_1 EN_RO_2_1 gnd 0
V_EN_RO_2_2 EN_RO_2_2 gnd 1
V_EN_RO_2_3 EN_RO_2_3 gnd 1
V_EN_RO_2_4 EN_RO_2_4 gnd 0
V_EN_RO_2_5 EN_RO_2_5 gnd 0
V_EN_RO_2_6 EN_RO_2_6 gnd 0
V_EN_RO_2_7 EN_RO_2_7 gnd 0
V_EN_RO_2_8 EN_RO_2_8 gnd 0
V_EN_RO_2_9 EN_RO_2_9 gnd 0
V_EN_RO_3_0 EN_RO_3_0 gnd 1
V_EN_RO_3_1 EN_RO_3_1 gnd 1
V_EN_RO_3_2 EN_RO_3_2 gnd 1
V_EN_RO_3_3 EN_RO_3_3 gnd 0
V_EN_RO_3_4 EN_RO_3_4 gnd 0
V_EN_RO_3_5 EN_RO_3_5 gnd 1
V_EN_RO_3_6 EN_RO_3_6 gnd 1
V_EN_RO_3_7 EN_RO_3_7 gnd 0
V_EN_RO_3_8 EN_RO_3_8 gnd 1
V_EN_RO_3_9 EN_RO_3_9 gnd 0
V_EN_RO_4_0 EN_RO_4_0 gnd 1
V_EN_RO_4_1 EN_RO_4_1 gnd 1
V_EN_RO_4_2 EN_RO_4_2 gnd 1
V_EN_RO_4_3 EN_RO_4_3 gnd 1
V_EN_RO_4_4 EN_RO_4_4 gnd 0
V_EN_RO_4_5 EN_RO_4_5 gnd 0
V_EN_RO_4_6 EN_RO_4_6 gnd 0
V_EN_RO_4_7 EN_RO_4_7 gnd 1
V_EN_RO_4_8 EN_RO_4_8 gnd 1
V_EN_RO_4_9 EN_RO_4_9 gnd 1
V_EN_RO_5_0 EN_RO_5_0 gnd 1
V_EN_RO_5_1 EN_RO_5_1 gnd 1
V_EN_RO_5_2 EN_RO_5_2 gnd 1
V_EN_RO_5_3 EN_RO_5_3 gnd 0
V_EN_RO_5_4 EN_RO_5_4 gnd 1
V_EN_RO_5_5 EN_RO_5_5 gnd 1
V_EN_RO_5_6 EN_RO_5_6 gnd 1
V_EN_RO_5_7 EN_RO_5_7 gnd 0
V_EN_RO_5_8 EN_RO_5_8 gnd 1
V_EN_RO_5_9 EN_RO_5_9 gnd 0
V_EN_RO_6_0 EN_RO_6_0 gnd 0
V_EN_RO_6_1 EN_RO_6_1 gnd 1
V_EN_RO_6_2 EN_RO_6_2 gnd 1
V_EN_RO_6_3 EN_RO_6_3 gnd 0
V_EN_RO_6_4 EN_RO_6_4 gnd 1
V_EN_RO_6_5 EN_RO_6_5 gnd 0
V_EN_RO_6_6 EN_RO_6_6 gnd 1
V_EN_RO_6_7 EN_RO_6_7 gnd 0
V_EN_RO_6_8 EN_RO_6_8 gnd 0
V_EN_RO_6_9 EN_RO_6_9 gnd 0
V_EN_RO_7_0 EN_RO_7_0 gnd 1
V_EN_RO_7_1 EN_RO_7_1 gnd 1
V_EN_RO_7_2 EN_RO_7_2 gnd 0
V_EN_RO_7_3 EN_RO_7_3 gnd 0
V_EN_RO_7_4 EN_RO_7_4 gnd 0
V_EN_RO_7_5 EN_RO_7_5 gnd 1
V_EN_RO_7_6 EN_RO_7_6 gnd 1
V_EN_RO_7_7 EN_RO_7_7 gnd 0
V_EN_RO_7_8 EN_RO_7_8 gnd 0
V_EN_RO_7_9 EN_RO_7_9 gnd 1
V_EN_RO_8_0 EN_RO_8_0 gnd 1
V_EN_RO_8_1 EN_RO_8_1 gnd 0
V_EN_RO_8_2 EN_RO_8_2 gnd 0
V_EN_RO_8_3 EN_RO_8_3 gnd 1
V_EN_RO_8_4 EN_RO_8_4 gnd 0
V_EN_RO_8_5 EN_RO_8_5 gnd 1
V_EN_RO_8_6 EN_RO_8_6 gnd 0
V_EN_RO_8_7 EN_RO_8_7 gnd 0
V_EN_RO_8_8 EN_RO_8_8 gnd 1
V_EN_RO_8_9 EN_RO_8_9 gnd 0
V_EN_RO_9_0 EN_RO_9_0 gnd 0
V_EN_RO_9_1 EN_RO_9_1 gnd 1
V_EN_RO_9_2 EN_RO_9_2 gnd 1
V_EN_RO_9_3 EN_RO_9_3 gnd 0
V_EN_RO_9_4 EN_RO_9_4 gnd 1
V_EN_RO_9_5 EN_RO_9_5 gnd 0
V_EN_RO_9_6 EN_RO_9_6 gnd 1
V_EN_RO_9_7 EN_RO_9_7 gnd 1
V_EN_RO_9_8 EN_RO_9_8 gnd 1
V_EN_RO_9_9 EN_RO_9_9 gnd 0

* Coupler enables
V_EN_C_0_0__0_1 EN_C_0_0__0_1 gnd 0
V_EN_C_0_0__1_0 EN_C_0_0__1_0 gnd 1
V_EN_C_0_1__0_2 EN_C_0_1__0_2 gnd 0
V_EN_C_0_1__1_0 EN_C_0_1__1_0 gnd 0
V_EN_C_0_1__1_1 EN_C_0_1__1_1 gnd 0
V_EN_C_0_2__0_3 EN_C_0_2__0_3 gnd 0
V_EN_C_0_2__1_1 EN_C_0_2__1_1 gnd 0
V_EN_C_0_2__1_2 EN_C_0_2__1_2 gnd 0
V_EN_C_0_3__0_4 EN_C_0_3__0_4 gnd 0
V_EN_C_0_3__1_2 EN_C_0_3__1_2 gnd 0
V_EN_C_0_3__1_3 EN_C_0_3__1_3 gnd 0
V_EN_C_0_4__0_5 EN_C_0_4__0_5 gnd 0
V_EN_C_0_4__1_3 EN_C_0_4__1_3 gnd 0
V_EN_C_0_4__1_4 EN_C_0_4__1_4 gnd 0
V_EN_C_0_5__0_6 EN_C_0_5__0_6 gnd 0
V_EN_C_0_5__1_4 EN_C_0_5__1_4 gnd 0
V_EN_C_0_5__1_5 EN_C_0_5__1_5 gnd 0
V_EN_C_0_6__0_7 EN_C_0_6__0_7 gnd 0
V_EN_C_0_6__1_5 EN_C_0_6__1_5 gnd 0
V_EN_C_0_6__1_6 EN_C_0_6__1_6 gnd 0
V_EN_C_0_7__0_8 EN_C_0_7__0_8 gnd 1
V_EN_C_0_7__1_6 EN_C_0_7__1_6 gnd 0
V_EN_C_0_7__1_7 EN_C_0_7__1_7 gnd 0
V_EN_C_0_8__0_9 EN_C_0_8__0_9 gnd 0
V_EN_C_0_8__1_7 EN_C_0_8__1_7 gnd 0
V_EN_C_0_8__1_8 EN_C_0_8__1_8 gnd 0
V_EN_C_0_9__1_8 EN_C_0_9__1_8 gnd 0
V_EN_C_0_9__1_9 EN_C_0_9__1_9 gnd 0
V_EN_C_1_0__1_1 EN_C_1_0__1_1 gnd 0
V_EN_C_1_0__2_0 EN_C_1_0__2_0 gnd 1
V_EN_C_1_0__2_1 EN_C_1_0__2_1 gnd 0
V_EN_C_1_1__1_2 EN_C_1_1__1_2 gnd 0
V_EN_C_1_1__2_1 EN_C_1_1__2_1 gnd 0
V_EN_C_1_1__2_2 EN_C_1_1__2_2 gnd 0
V_EN_C_1_2__1_3 EN_C_1_2__1_3 gnd 0
V_EN_C_1_2__2_2 EN_C_1_2__2_2 gnd 0
V_EN_C_1_2__2_3 EN_C_1_2__2_3 gnd 0
V_EN_C_1_3__1_4 EN_C_1_3__1_4 gnd 1
V_EN_C_1_3__2_3 EN_C_1_3__2_3 gnd 1
V_EN_C_1_3__2_4 EN_C_1_3__2_4 gnd 0
V_EN_C_1_4__1_5 EN_C_1_4__1_5 gnd 1
V_EN_C_1_4__2_4 EN_C_1_4__2_4 gnd 0
V_EN_C_1_4__2_5 EN_C_1_4__2_5 gnd 0
V_EN_C_1_5__1_6 EN_C_1_5__1_6 gnd 0
V_EN_C_1_5__2_5 EN_C_1_5__2_5 gnd 0
V_EN_C_1_5__2_6 EN_C_1_5__2_6 gnd 0
V_EN_C_1_6__1_7 EN_C_1_6__1_7 gnd 0
V_EN_C_1_6__2_6 EN_C_1_6__2_6 gnd 0
V_EN_C_1_6__2_7 EN_C_1_6__2_7 gnd 0
V_EN_C_1_7__1_8 EN_C_1_7__1_8 gnd 0
V_EN_C_1_7__2_7 EN_C_1_7__2_7 gnd 0
V_EN_C_1_7__2_8 EN_C_1_7__2_8 gnd 0
V_EN_C_1_8__1_9 EN_C_1_8__1_9 gnd 0
V_EN_C_1_8__2_8 EN_C_1_8__2_8 gnd 0
V_EN_C_1_8__2_9 EN_C_1_8__2_9 gnd 0
V_EN_C_1_9__2_9 EN_C_1_9__2_9 gnd 0
V_EN_C_2_0__2_1 EN_C_2_0__2_1 gnd 0
V_EN_C_2_0__3_0 EN_C_2_0__3_0 gnd 1
V_EN_C_2_1__2_2 EN_C_2_1__2_2 gnd 0
V_EN_C_2_1__3_0 EN_C_2_1__3_0 gnd 0
V_EN_C_2_1__3_1 EN_C_2_1__3_1 gnd 0
V_EN_C_2_2__2_3 EN_C_2_2__2_3 gnd 1
V_EN_C_2_2__3_1 EN_C_2_2__3_1 gnd 0
V_EN_C_2_2__3_2 EN_C_2_2__3_2 gnd 1
V_EN_C_2_3__2_4 EN_C_2_3__2_4 gnd 0
V_EN_C_2_3__3_2 EN_C_2_3__3_2 gnd 1
V_EN_C_2_3__3_3 EN_C_2_3__3_3 gnd 0
V_EN_C_2_4__2_5 EN_C_2_4__2_5 gnd 0
V_EN_C_2_4__3_3 EN_C_2_4__3_3 gnd 0
V_EN_C_2_4__3_4 EN_C_2_4__3_4 gnd 0
V_EN_C_2_5__2_6 EN_C_2_5__2_6 gnd 0
V_EN_C_2_5__3_4 EN_C_2_5__3_4 gnd 0
V_EN_C_2_5__3_5 EN_C_2_5__3_5 gnd 0
V_EN_C_2_6__2_7 EN_C_2_6__2_7 gnd 0
V_EN_C_2_6__3_5 EN_C_2_6__3_5 gnd 0
V_EN_C_2_6__3_6 EN_C_2_6__3_6 gnd 0
V_EN_C_2_7__2_8 EN_C_2_7__2_8 gnd 0
V_EN_C_2_7__3_6 EN_C_2_7__3_6 gnd 0
V_EN_C_2_7__3_7 EN_C_2_7__3_7 gnd 0
V_EN_C_2_8__2_9 EN_C_2_8__2_9 gnd 0
V_EN_C_2_8__3_7 EN_C_2_8__3_7 gnd 0
V_EN_C_2_8__3_8 EN_C_2_8__3_8 gnd 0
V_EN_C_2_9__3_8 EN_C_2_9__3_8 gnd 0
V_EN_C_2_9__3_9 EN_C_2_9__3_9 gnd 0
V_EN_C_3_0__3_1 EN_C_3_0__3_1 gnd 1
V_EN_C_3_0__4_0 EN_C_3_0__4_0 gnd 0
V_EN_C_3_0__4_1 EN_C_3_0__4_1 gnd 0
V_EN_C_3_1__3_2 EN_C_3_1__3_2 gnd 1
V_EN_C_3_1__4_1 EN_C_3_1__4_1 gnd 1
V_EN_C_3_1__4_2 EN_C_3_1__4_2 gnd 0
V_EN_C_3_2__3_3 EN_C_3_2__3_3 gnd 0
V_EN_C_3_2__4_2 EN_C_3_2__4_2 gnd 1
V_EN_C_3_2__4_3 EN_C_3_2__4_3 gnd 1
V_EN_C_3_3__3_4 EN_C_3_3__3_4 gnd 0
V_EN_C_3_3__4_3 EN_C_3_3__4_3 gnd 0
V_EN_C_3_3__4_4 EN_C_3_3__4_4 gnd 0
V_EN_C_3_4__3_5 EN_C_3_4__3_5 gnd 0
V_EN_C_3_4__4_4 EN_C_3_4__4_4 gnd 0
V_EN_C_3_4__4_5 EN_C_3_4__4_5 gnd 0
V_EN_C_3_5__3_6 EN_C_3_5__3_6 gnd 1
V_EN_C_3_5__4_5 EN_C_3_5__4_5 gnd 0
V_EN_C_3_5__4_6 EN_C_3_5__4_6 gnd 0
V_EN_C_3_6__3_7 EN_C_3_6__3_7 gnd 0
V_EN_C_3_6__4_6 EN_C_3_6__4_6 gnd 0
V_EN_C_3_6__4_7 EN_C_3_6__4_7 gnd 1
V_EN_C_3_7__3_8 EN_C_3_7__3_8 gnd 0
V_EN_C_3_7__4_7 EN_C_3_7__4_7 gnd 0
V_EN_C_3_7__4_8 EN_C_3_7__4_8 gnd 0
V_EN_C_3_8__3_9 EN_C_3_8__3_9 gnd 0
V_EN_C_3_8__4_8 EN_C_3_8__4_8 gnd 1
V_EN_C_3_8__4_9 EN_C_3_8__4_9 gnd 0
V_EN_C_3_9__4_9 EN_C_3_9__4_9 gnd 0
V_EN_C_4_0__4_1 EN_C_4_0__4_1 gnd 1
V_EN_C_4_0__5_0 EN_C_4_0__5_0 gnd 0
V_EN_C_4_1__4_2 EN_C_4_1__4_2 gnd 1
V_EN_C_4_1__5_0 EN_C_4_1__5_0 gnd 1
V_EN_C_4_1__5_1 EN_C_4_1__5_1 gnd 1
V_EN_C_4_2__4_3 EN_C_4_2__4_3 gnd 0
V_EN_C_4_2__5_1 EN_C_4_2__5_1 gnd 1
V_EN_C_4_2__5_2 EN_C_4_2__5_2 gnd 1
V_EN_C_4_3__4_4 EN_C_4_3__4_4 gnd 0
V_EN_C_4_3__5_2 EN_C_4_3__5_2 gnd 0
V_EN_C_4_3__5_3 EN_C_4_3__5_3 gnd 0
V_EN_C_4_4__4_5 EN_C_4_4__4_5 gnd 0
V_EN_C_4_4__5_3 EN_C_4_4__5_3 gnd 0
V_EN_C_4_4__5_4 EN_C_4_4__5_4 gnd 0
V_EN_C_4_5__4_6 EN_C_4_5__4_6 gnd 0
V_EN_C_4_5__5_4 EN_C_4_5__5_4 gnd 0
V_EN_C_4_5__5_5 EN_C_4_5__5_5 gnd 0
V_EN_C_4_6__4_7 EN_C_4_6__4_7 gnd 0
V_EN_C_4_6__5_5 EN_C_4_6__5_5 gnd 0
V_EN_C_4_6__5_6 EN_C_4_6__5_6 gnd 0
V_EN_C_4_7__4_8 EN_C_4_7__4_8 gnd 1
V_EN_C_4_7__5_6 EN_C_4_7__5_6 gnd 1
V_EN_C_4_7__5_7 EN_C_4_7__5_7 gnd 0
V_EN_C_4_8__4_9 EN_C_4_8__4_9 gnd 1
V_EN_C_4_8__5_7 EN_C_4_8__5_7 gnd 0
V_EN_C_4_8__5_8 EN_C_4_8__5_8 gnd 1
V_EN_C_4_9__5_8 EN_C_4_9__5_8 gnd 1
V_EN_C_4_9__5_9 EN_C_4_9__5_9 gnd 0
V_EN_C_5_0__5_1 EN_C_5_0__5_1 gnd 1
V_EN_C_5_0__6_0 EN_C_5_0__6_0 gnd 0
V_EN_C_5_0__6_1 EN_C_5_0__6_1 gnd 1
V_EN_C_5_1__5_2 EN_C_5_1__5_2 gnd 0
V_EN_C_5_1__6_1 EN_C_5_1__6_1 gnd 1
V_EN_C_5_1__6_2 EN_C_5_1__6_2 gnd 1
V_EN_C_5_2__5_3 EN_C_5_2__5_3 gnd 0
V_EN_C_5_2__6_2 EN_C_5_2__6_2 gnd 0
V_EN_C_5_2__6_3 EN_C_5_2__6_3 gnd 0
V_EN_C_5_3__5_4 EN_C_5_3__5_4 gnd 0
V_EN_C_5_3__6_3 EN_C_5_3__6_3 gnd 0
V_EN_C_5_3__6_4 EN_C_5_3__6_4 gnd 0
V_EN_C_5_4__5_5 EN_C_5_4__5_5 gnd 1
V_EN_C_5_4__6_4 EN_C_5_4__6_4 gnd 1
V_EN_C_5_4__6_5 EN_C_5_4__6_5 gnd 0
V_EN_C_5_5__5_6 EN_C_5_5__5_6 gnd 1
V_EN_C_5_5__6_5 EN_C_5_5__6_5 gnd 0
V_EN_C_5_5__6_6 EN_C_5_5__6_6 gnd 1
V_EN_C_5_6__5_7 EN_C_5_6__5_7 gnd 0
V_EN_C_5_6__6_6 EN_C_5_6__6_6 gnd 1
V_EN_C_5_6__6_7 EN_C_5_6__6_7 gnd 0
V_EN_C_5_7__5_8 EN_C_5_7__5_8 gnd 0
V_EN_C_5_7__6_7 EN_C_5_7__6_7 gnd 0
V_EN_C_5_7__6_8 EN_C_5_7__6_8 gnd 0
V_EN_C_5_8__5_9 EN_C_5_8__5_9 gnd 0
V_EN_C_5_8__6_8 EN_C_5_8__6_8 gnd 0
V_EN_C_5_8__6_9 EN_C_5_8__6_9 gnd 0
V_EN_C_5_9__6_9 EN_C_5_9__6_9 gnd 0
V_EN_C_6_0__6_1 EN_C_6_0__6_1 gnd 0
V_EN_C_6_0__7_0 EN_C_6_0__7_0 gnd 0
V_EN_C_6_1__6_2 EN_C_6_1__6_2 gnd 1
V_EN_C_6_1__7_0 EN_C_6_1__7_0 gnd 1
V_EN_C_6_1__7_1 EN_C_6_1__7_1 gnd 1
V_EN_C_6_2__6_3 EN_C_6_2__6_3 gnd 0
V_EN_C_6_2__7_1 EN_C_6_2__7_1 gnd 0
V_EN_C_6_2__7_2 EN_C_6_2__7_2 gnd 0
V_EN_C_6_3__6_4 EN_C_6_3__6_4 gnd 0
V_EN_C_6_3__7_2 EN_C_6_3__7_2 gnd 0
V_EN_C_6_3__7_3 EN_C_6_3__7_3 gnd 0
V_EN_C_6_4__6_5 EN_C_6_4__6_5 gnd 0
V_EN_C_6_4__7_3 EN_C_6_4__7_3 gnd 0
V_EN_C_6_4__7_4 EN_C_6_4__7_4 gnd 0
V_EN_C_6_5__6_6 EN_C_6_5__6_6 gnd 0
V_EN_C_6_5__7_4 EN_C_6_5__7_4 gnd 0
V_EN_C_6_5__7_5 EN_C_6_5__7_5 gnd 0
V_EN_C_6_6__6_7 EN_C_6_6__6_7 gnd 0
V_EN_C_6_6__7_5 EN_C_6_6__7_5 gnd 1
V_EN_C_6_6__7_6 EN_C_6_6__7_6 gnd 1
V_EN_C_6_7__6_8 EN_C_6_7__6_8 gnd 0
V_EN_C_6_7__7_6 EN_C_6_7__7_6 gnd 0
V_EN_C_6_7__7_7 EN_C_6_7__7_7 gnd 0
V_EN_C_6_8__6_9 EN_C_6_8__6_9 gnd 0
V_EN_C_6_8__7_7 EN_C_6_8__7_7 gnd 0
V_EN_C_6_8__7_8 EN_C_6_8__7_8 gnd 0
V_EN_C_6_9__7_8 EN_C_6_9__7_8 gnd 0
V_EN_C_6_9__7_9 EN_C_6_9__7_9 gnd 0
V_EN_C_7_0__7_1 EN_C_7_0__7_1 gnd 0
V_EN_C_7_0__8_0 EN_C_7_0__8_0 gnd 1
V_EN_C_7_0__8_1 EN_C_7_0__8_1 gnd 0
V_EN_C_7_1__7_2 EN_C_7_1__7_2 gnd 0
V_EN_C_7_1__8_1 EN_C_7_1__8_1 gnd 0
V_EN_C_7_1__8_2 EN_C_7_1__8_2 gnd 0
V_EN_C_7_2__7_3 EN_C_7_2__7_3 gnd 0
V_EN_C_7_2__8_2 EN_C_7_2__8_2 gnd 0
V_EN_C_7_2__8_3 EN_C_7_2__8_3 gnd 0
V_EN_C_7_3__7_4 EN_C_7_3__7_4 gnd 0
V_EN_C_7_3__8_3 EN_C_7_3__8_3 gnd 0
V_EN_C_7_3__8_4 EN_C_7_3__8_4 gnd 0
V_EN_C_7_4__7_5 EN_C_7_4__7_5 gnd 0
V_EN_C_7_4__8_4 EN_C_7_4__8_4 gnd 0
V_EN_C_7_4__8_5 EN_C_7_4__8_5 gnd 0
V_EN_C_7_5__7_6 EN_C_7_5__7_6 gnd 0
V_EN_C_7_5__8_5 EN_C_7_5__8_5 gnd 1
V_EN_C_7_5__8_6 EN_C_7_5__8_6 gnd 0
V_EN_C_7_6__7_7 EN_C_7_6__7_7 gnd 0
V_EN_C_7_6__8_6 EN_C_7_6__8_6 gnd 0
V_EN_C_7_6__8_7 EN_C_7_6__8_7 gnd 0
V_EN_C_7_7__7_8 EN_C_7_7__7_8 gnd 0
V_EN_C_7_7__8_7 EN_C_7_7__8_7 gnd 0
V_EN_C_7_7__8_8 EN_C_7_7__8_8 gnd 0
V_EN_C_7_8__7_9 EN_C_7_8__7_9 gnd 0
V_EN_C_7_8__8_8 EN_C_7_8__8_8 gnd 0
V_EN_C_7_8__8_9 EN_C_7_8__8_9 gnd 0
V_EN_C_7_9__8_9 EN_C_7_9__8_9 gnd 0
V_EN_C_8_0__8_1 EN_C_8_0__8_1 gnd 0
V_EN_C_8_0__9_0 EN_C_8_0__9_0 gnd 0
V_EN_C_8_1__8_2 EN_C_8_1__8_2 gnd 0
V_EN_C_8_1__9_0 EN_C_8_1__9_0 gnd 0
V_EN_C_8_1__9_1 EN_C_8_1__9_1 gnd 0
V_EN_C_8_2__8_3 EN_C_8_2__8_3 gnd 0
V_EN_C_8_2__9_1 EN_C_8_2__9_1 gnd 0
V_EN_C_8_2__9_2 EN_C_8_2__9_2 gnd 0
V_EN_C_8_3__8_4 EN_C_8_3__8_4 gnd 0
V_EN_C_8_3__9_2 EN_C_8_3__9_2 gnd 1
V_EN_C_8_3__9_3 EN_C_8_3__9_3 gnd 0
V_EN_C_8_4__8_5 EN_C_8_4__8_5 gnd 0
V_EN_C_8_4__9_3 EN_C_8_4__9_3 gnd 0
V_EN_C_8_4__9_4 EN_C_8_4__9_4 gnd 0
V_EN_C_8_5__8_6 EN_C_8_5__8_6 gnd 0
V_EN_C_8_5__9_4 EN_C_8_5__9_4 gnd 1
V_EN_C_8_5__9_5 EN_C_8_5__9_5 gnd 0
V_EN_C_8_6__8_7 EN_C_8_6__8_7 gnd 0
V_EN_C_8_6__9_5 EN_C_8_6__9_5 gnd 0
V_EN_C_8_6__9_6 EN_C_8_6__9_6 gnd 0
V_EN_C_8_7__8_8 EN_C_8_7__8_8 gnd 0
V_EN_C_8_7__9_6 EN_C_8_7__9_6 gnd 0
V_EN_C_8_7__9_7 EN_C_8_7__9_7 gnd 0
V_EN_C_8_8__8_9 EN_C_8_8__8_9 gnd 0
V_EN_C_8_8__9_7 EN_C_8_8__9_7 gnd 1
V_EN_C_8_8__9_8 EN_C_8_8__9_8 gnd 1
V_EN_C_8_9__9_8 EN_C_8_9__9_8 gnd 0
V_EN_C_8_9__9_9 EN_C_8_9__9_9 gnd 0
V_EN_C_9_0__9_1 EN_C_9_0__9_1 gnd 0
V_EN_C_9_1__9_2 EN_C_9_1__9_2 gnd 1
V_EN_C_9_2__9_3 EN_C_9_2__9_3 gnd 0
V_EN_C_9_3__9_4 EN_C_9_3__9_4 gnd 0
V_EN_C_9_4__9_5 EN_C_9_4__9_5 gnd 0
V_EN_C_9_5__9_6 EN_C_9_5__9_6 gnd 0
V_EN_C_9_6__9_7 EN_C_9_6__9_7 gnd 1
V_EN_C_9_7__9_8 EN_C_9_7__9_8 gnd 1
V_EN_C_9_8__9_9 EN_C_9_8__9_9 gnd 0

VDD vdd gnd 1.0

.control
save time N_0_0_1 N_0_1_1 N_0_2_1 N_0_3_1 N_0_4_1 N_0_5_1 N_0_6_1 N_0_7_1 N_0_8_1 N_0_9_1 N_1_0_1 N_1_1_1 N_1_2_1 N_1_3_1 N_1_4_1 N_1_5_1 N_1_6_1 N_1_7_1 N_1_8_1 N_1_9_1 N_2_0_1 N_2_1_1 N_2_2_1 N_2_3_1 N_2_4_1 N_2_5_1 N_2_6_1 N_2_7_1 N_2_8_1 N_2_9_1 N_3_0_1 N_3_1_1 N_3_2_1 N_3_3_1 N_3_4_1 N_3_5_1 N_3_6_1 N_3_7_1 N_3_8_1 N_3_9_1 N_4_0_1 N_4_1_1 N_4_2_1 N_4_3_1 N_4_4_1 N_4_5_1 N_4_6_1 N_4_7_1 N_4_8_1 N_4_9_1 N_5_0_1 N_5_1_1 N_5_2_1 N_5_3_1 N_5_4_1 N_5_5_1 N_5_6_1 N_5_7_1 N_5_8_1 N_5_9_1 N_6_0_1 N_6_1_1 N_6_2_1 N_6_3_1 N_6_4_1 N_6_5_1 N_6_6_1 N_6_7_1 N_6_8_1 N_6_9_1 N_7_0_1 N_7_1_1 N_7_2_1 N_7_3_1 N_7_4_1 N_7_5_1 N_7_6_1 N_7_7_1 N_7_8_1 N_7_9_1 N_8_0_1 N_8_1_1 N_8_2_1 N_8_3_1 N_8_4_1 N_8_5_1 N_8_6_1 N_8_7_1 N_8_8_1 N_8_9_1 N_9_0_1 N_9_1_1 N_9_2_1 N_9_3_1 N_9_4_1 N_9_5_1 N_9_6_1 N_9_7_1 N_9_8_1 N_9_9_1
tran 0.1ns 2us uic
set filetype=ascii
set wr_singlescale
set wr_vecnames
set csvdelim=comma
wrdata output_nodes.csv time N_0_0_1 N_0_1_1 N_0_2_1 N_0_3_1 N_0_4_1 N_0_5_1 N_0_6_1 N_0_7_1 N_0_8_1 N_0_9_1 N_1_0_1 N_1_1_1 N_1_2_1 N_1_3_1 N_1_4_1 N_1_5_1 N_1_6_1 N_1_7_1 N_1_8_1 N_1_9_1 N_2_0_1 N_2_1_1 N_2_2_1 N_2_3_1 N_2_4_1 N_2_5_1 N_2_6_1 N_2_7_1 N_2_8_1 N_2_9_1 N_3_0_1 N_3_1_1 N_3_2_1 N_3_3_1 N_3_4_1 N_3_5_1 N_3_6_1 N_3_7_1 N_3_8_1 N_3_9_1 N_4_0_1 N_4_1_1 N_4_2_1 N_4_3_1 N_4_4_1 N_4_5_1 N_4_6_1 N_4_7_1 N_4_8_1 N_4_9_1 N_5_0_1 N_5_1_1 N_5_2_1 N_5_3_1 N_5_4_1 N_5_5_1 N_5_6_1 N_5_7_1 N_5_8_1 N_5_9_1 N_6_0_1 N_6_1_1 N_6_2_1 N_6_3_1 N_6_4_1 N_6_5_1 N_6_6_1 N_6_7_1 N_6_8_1 N_6_9_1 N_7_0_1 N_7_1_1 N_7_2_1 N_7_3_1 N_7_4_1 N_7_5_1 N_7_6_1 N_7_7_1 N_7_8_1 N_7_9_1 N_8_0_1 N_8_1_1 N_8_2_1 N_8_3_1 N_8_4_1 N_8_5_1 N_8_6_1 N_8_7_1 N_8_8_1 N_8_9_1 N_9_0_1 N_9_1_1 N_9_2_1 N_9_3_1 N_9_4_1 N_9_5_1 N_9_6_1 N_9_7_1 N_9_8_1 N_9_9_1
quit
.endc

.end
